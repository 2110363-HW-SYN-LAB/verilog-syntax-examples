// alternative syntax easier to read and beautiful code

module better_and_gate (
    input  wire a,
    input  wire b,
    output wire out
);

    assign out = a & b;

endmodule
