// alternative syntax easier to read and beautiful code

module better_and_gate (
    input  a,
    input  b,
    output out
);

    assign out = a & b;

endmodule
